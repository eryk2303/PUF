

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package sha256_typ is


		type function_initial_values is array(0 to 7) of std_logic_vector(31 downto 0);
		type constants_value_sha256 is array(0 to 63) of std_logic_vector(31 downto 0);


end sha256_typ;

package body sha256_typ is

end sha256_typ;
